LIBRARY IEEE;
USE IEEE.std_Logic_1164.all;
USE IEEE.Numeric_std.all;

--------------------------------------------------------------------------------
--                                                                            --
-- Global Parameters - values governed by external requirements               --
--                                                                            --
--------------------------------------------------------------------------------

PACKAGE fib_parameters IS
    CONSTANT BusWidth : INTEGER := 8;
END fib_parameters;
  
PACKAGE BODY fib_parameters IS
END PACKAGE BODY fib_parameters;