LIBRARY IEEE;
USE IEEE.Std_Logic_1164.ALL;
USE IEEE.Numeric_Std.ALL;

--------------------------------------------------------------------------------
--                                                                            --
-- Global Parameters - values governed by external requirements               --
--                                                                            --
--------------------------------------------------------------------------------

PACKAGE fib_parameters IS
    CONSTANT BusWidth : INTEGER := 8;
END fib_parameters;
  
PACKAGE BODY fib_parameters IS
END PACKAGE BODY fib_parameters;