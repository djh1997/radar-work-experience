LIBRARY IEEE;
USE IEEE.std_Logic_1164.ALL;
USE IEEE.Numeric_std.ALL;

--------------------------------------------------------------------------------
--                                                                            --
-- Global Parameters - values governed by external requirements               --
--                                                                            --
--------------------------------------------------------------------------------

PACKAGE fib_parameters IS
  CONSTANT BusWidth : INTEGER := 8;
END fib_parameters;

PACKAGE BODY fib_parameters IS
END PACKAGE BODY fib_parameters;